package afifo_test_pkg;
  import afifo_pkg::*;
  import afifo_rd_agent_pkg::*;
  import afifo_wr_agent_pkg::*;
  import afifo_env_pkg::*;
  import afifo_seq_pkg::*;
  `include "afifo_test_base.sv"
endpackage

package afifo_rd_agent_pkg;
  import afifo_pkg::*;
  `include "afifo_rd_txn.svh"
  `include "afifo_rd_driver.svh"
  `include "afifo_rd_monitor.svh"
  `include "afifo_rd_agent.svh"
endpackage

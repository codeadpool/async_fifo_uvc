`ifndef AFIFO_WR_PKG
`define AFIFO_WR_PKG
package afifo_wr_pkg;
  import uvm_pkg::*; 
  `include "uvm_macros.svh"


endpackage
`endif

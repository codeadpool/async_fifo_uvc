package afifo_tb_pkg;
  import afifo_pkg::*;
  import afifo_rd_agent_pkg::*;
  import afifo_wr_agent_pkg::*;
  import afifo_env_pkg::*;
  import afifo_seq_pkg::*;
  import afifo_test_pkg::*;
  import tb_params_pkg::*;
endpackage

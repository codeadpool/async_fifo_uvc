package afifo_wr_agent_pkg;
  import afifo_pkg::*;
  `include "afifo_wr_txn.svh"
  `include "afifo_wr_driver.svh"
  `include "afifo_wr_monitor.svh"
  `include "afifo_wr_driver_bfm.svh"
  `include "afifo_wr_monitor_bfm.svh"

  `include "afifo_wr_agent.svh"
endpackage

package afifo_env_pkg;
  import afifo_pkg::*;
  import afifo_rd_agent_pkg::*;
  import afifo_wr_agent_pkg::*;
  `include "afifo_scoreboard.svh"
  `include "afifo_env.svh"
endpackage

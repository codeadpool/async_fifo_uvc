package afifo_pkg;
  `include "afifo_mcseqr.svh"
endpackage

package afifo_seq_pkg;
  import afifo_pkg::*;
  import afifo_rd_agent_pkg::*;
  import afifo_wr_agent_pkg::*;
  `include "afifo_seq_lib.svh"
  `include "afifo_vseq_lib.svh"
endpackage
